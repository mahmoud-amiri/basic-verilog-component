module moduleName #(
    parameter AND_OUTPUTS_WIDTH = 10
)
(
    input clk,
    input reset_n,
    output [AND_OUTPUTS_WIDTH-1:0] output,

);
    
endmodule
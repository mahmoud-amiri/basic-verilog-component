interface AndGateIf;
    logic a, b; // Inputs
    logic y;    // Output
endinterface

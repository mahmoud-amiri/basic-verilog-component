package pkg;

`include "driver.sv"
`include "interface.sv"
`include "coverage.sv"
//`include "firewall.sv"
`include "monitor.sv"
`include "scoreoard.sv"
`include "sequenceitem.sv"
`include "sequencer.sv"
`include "agent.sv"
`include "environment.sv"

endpackage : pkg